CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
48 106 1872 1004
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 106 1872 1004
143654930 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 761 649 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 773 598 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 762 451 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 766 416 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 283 243 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 281 321 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-7 -24 7 -16
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 307 276 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 290 180 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3747 0 0
0
0
9 2-In NOR~
219 1171 508 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3549 0 0
0
0
14 Logic Display~
6 1282 489 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
8 2-In OR~
219 911 618 0 3 22
0 5 6 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
9325 0 0
0
0
8 2-In OR~
219 1005 479 0 3 22
0 7 8 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
8903 0 0
0
0
9 Inverter~
13 839 548 0 2 22
0 10 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3834 0 0
0
0
9 2-In AND~
219 909 539 0 3 22
0 9 11 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3363 0 0
0
0
9 2-In AND~
219 907 429 0 3 22
0 10 9 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7668 0 0
0
0
14 Logic Display~
6 823 231 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4718 0 0
0
0
14 Logic Display~
6 737 233 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3874 0 0
0
0
8 2-In OR~
219 423 300 0 3 22
0 15 14 17
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6671 0 0
0
0
8 2-In OR~
219 417 230 0 3 22
0 16 13 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3789 0 0
0
0
9 2-In AND~
219 576 256 0 3 22
0 18 17 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4871 0 0
0
0
21
3 0 2 0 0 4096 0 9 0 0 2 2
1210 508
1210 507
0 1 2 0 0 8320 0 0 10 0 0 3
1205 508
1205 507
1282 507
2 3 3 0 0 8320 0 9 11 0 0 5
1158 517
1158 517
1029 517
1029 618
944 618
3 1 4 0 0 4224 0 12 9 0 0 5
1038 479
1145 479
1145 499
1158 499
1158 499
1 1 5 0 0 4224 0 2 11 0 0 4
785 598
899 598
899 609
898 609
1 2 6 0 0 4224 0 1 11 0 0 3
773 649
898 649
898 627
3 1 7 0 0 4224 0 15 12 0 0 4
928 429
986 429
986 470
992 470
3 2 8 0 0 4224 0 14 12 0 0 4
930 539
983 539
983 488
992 488
1 0 9 0 0 8192 0 14 0 0 11 3
885 530
856 530
856 438
0 1 10 0 0 4096 0 0 13 12 0 5
843 420
843 514
816 514
816 548
824 548
1 2 9 0 0 8320 0 3 15 0 0 3
774 451
774 438
883 438
1 1 10 0 0 8320 0 4 15 0 0 3
778 416
778 420
883 420
2 2 11 0 0 4224 0 13 14 0 0 2
860 548
885 548
1 1 12 0 0 8192 0 17 16 0 0 3
737 251
737 249
823 249
3 1 12 0 0 4224 0 20 17 0 0 3
597 256
737 256
737 251
1 2 13 0 0 4224 0 5 19 0 0 4
295 243
393 243
393 239
404 239
1 2 14 0 0 4224 0 6 18 0 0 4
293 321
398 321
398 309
410 309
1 1 15 0 0 4224 0 7 18 0 0 4
319 276
395 276
395 291
410 291
1 1 16 0 0 8320 0 8 19 0 0 3
302 180
302 221
404 221
3 2 17 0 0 4224 0 18 20 0 0 4
456 300
544 300
544 265
552 265
3 1 18 0 0 4224 0 19 20 0 0 4
450 230
544 230
544 247
552 247
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
712 632 728 656
722 640 730 656
1 d
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
708 584 724 608
718 592 726 608
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
719 392 735 416
726 399 734 415
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
715 434 731 458
725 442 733 458
1 b
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
